//==================================================================================================
//  Note:          Use only for teaching materials of IC Design Lab, NTHU.
//  Copyright: (c) 2022 Vision Circuits and Systems Lab, NTHU, Taiwan. ALL Rights Reserved.
//==================================================================================================


module enigma(clk, srst_n, load, encrypt, crypt_mode, table_idx, code_in, code_out, code_valid);
input clk;         // clock 
input srst_n;      // synchronous reset (active low)
input load;        // load control signal (level sensitive). 0/1: inactive/active
input encrypt;     // encrypt control signal (level sensitive). 0/1: inactive/active
input crypt_mode;  // 0: encrypt; 1:decrypt;
input [2-1:0] table_idx; // table_idx indicates which rotor to be loaded 
						             // 2'b00: rotorA
						             // 2'b01: rotorB
						             // 2'b10: plugboard
input [6-1:0] code_in;	// When load is active, then code_in is input of rotors. 
							          // When encrypy is active, then code_in is input of code words.
							          // Note: We only use rotorA in part1.
output reg [6-1:0] code_out;   // encrypted code word (register output)
output reg code_valid;         // 0: non-valid code_out; 1: valid code_out (register output)

reg load_buf;        
reg encrypt_buf;     
reg crypt_mode_buf;  
reg [1:0] table_idx_buf; 
reg [5:0] code_in_buf;
reg code_valid_nxt;
reg [5:0] rotorB_backward_pipe;
reg encrypt_pipe;

wire [5:0] rotorA [0:63];
wire [5:0] rotorB [0:63];
wire [5:0] plugboard [0:31];
wire [5:0] rotorA_forward;
wire [5:0] rotorB_forward;
wire [5:0] plugboard_forward;
wire [5:0] plugboard_backward;
wire [5:0] rotorB_backward;
wire [5:0] code_in_1;
wire [5:0] code_in_2;
wire [5:0] code_in_3;
wire [5:0] shift_accu; // shift rotorA
wire [5:0] shift_accu_pipe;
wire [5:0] shift_backward;
wire [5:0] rotorB_mode [0:63];
wire [5:0] code_out_nxt;

// sequential
always@(posedge clk) begin
    if(~srst_n) code_valid <= 0;
    else code_valid <= code_valid_nxt;
	load_buf <= load;
	encrypt_buf <= encrypt;
	crypt_mode_buf <= crypt_mode;
	table_idx_buf <= table_idx;
	code_in_buf <= code_in;
    code_out <= code_out_nxt;
    rotorB_backward_pipe <= rotorB_backward;
    encrypt_pipe <= encrypt_buf;
end

// other regs and signals
always @(*) code_valid_nxt = (encrypt_pipe) ? 1'b1 : 1'b0;


rotorA a(
	.clk(clk),
	.table_idx_buf(table_idx_buf),
	.load_buf(load_buf),
	.code_in_buf(code_in_buf),
	.shift_accu(shift_accu),
    .shift_backward(shift_backward),
	.rotorA0(rotorA[0]),
    .rotorA1(rotorA[1]),
    .rotorA2(rotorA[2]),
    .rotorA3(rotorA[3]),
    .rotorA4(rotorA[4]),
    .rotorA5(rotorA[5]),
    .rotorA6(rotorA[6]),
    .rotorA7(rotorA[7]),
    .rotorA8(rotorA[8]),
    .rotorA9(rotorA[9]),
    .rotorA10(rotorA[10]),
    .rotorA11(rotorA[11]),
    .rotorA12(rotorA[12]),
    .rotorA13(rotorA[13]),
    .rotorA14(rotorA[14]),
    .rotorA15(rotorA[15]),
    .rotorA16(rotorA[16]),
    .rotorA17(rotorA[17]),
    .rotorA18(rotorA[18]),
    .rotorA19(rotorA[19]),
    .rotorA20(rotorA[20]),
    .rotorA21(rotorA[21]),
    .rotorA22(rotorA[22]),
    .rotorA23(rotorA[23]),
    .rotorA24(rotorA[24]),
    .rotorA25(rotorA[25]),
    .rotorA26(rotorA[26]),
    .rotorA27(rotorA[27]),
    .rotorA28(rotorA[28]),
    .rotorA29(rotorA[29]),
    .rotorA30(rotorA[30]),
    .rotorA31(rotorA[31]),
    .rotorA32(rotorA[32]),
    .rotorA33(rotorA[33]),
    .rotorA34(rotorA[34]),
    .rotorA35(rotorA[35]),
    .rotorA36(rotorA[36]),
    .rotorA37(rotorA[37]),
    .rotorA38(rotorA[38]),
    .rotorA39(rotorA[39]),
    .rotorA40(rotorA[40]),
    .rotorA41(rotorA[41]),
    .rotorA42(rotorA[42]),
    .rotorA43(rotorA[43]),
    .rotorA44(rotorA[44]),
    .rotorA45(rotorA[45]),
    .rotorA46(rotorA[46]),
    .rotorA47(rotorA[47]),
    .rotorA48(rotorA[48]),
    .rotorA49(rotorA[49]),
    .rotorA50(rotorA[50]),
    .rotorA51(rotorA[51]),
    .rotorA52(rotorA[52]),
    .rotorA53(rotorA[53]),
    .rotorA54(rotorA[54]),
    .rotorA55(rotorA[55]),
    .rotorA56(rotorA[56]),
    .rotorA57(rotorA[57]),
    .rotorA58(rotorA[58]),
    .rotorA59(rotorA[59]),
    .rotorA60(rotorA[60]),
    .rotorA61(rotorA[61]),
    .rotorA62(rotorA[62]),
    .rotorA63(rotorA[63]),
	.code_in_1(code_in_1),
	.code_in_2(code_in_2),
	.code_in_3(code_in_3)
);

rotorB b(
	.clk(clk),
    .table_idx_buf(table_idx_buf),
    .load_buf(load_buf),
	.code_in_buf(code_in_buf),
	.rotorB_nxt0(rotorB_mode[0]),
    .rotorB_nxt1(rotorB_mode[1]),
    .rotorB_nxt2(rotorB_mode[2]),
    .rotorB_nxt3(rotorB_mode[3]),
    .rotorB_nxt4(rotorB_mode[4]),
    .rotorB_nxt5(rotorB_mode[5]),
    .rotorB_nxt6(rotorB_mode[6]),
    .rotorB_nxt7(rotorB_mode[7]),
    .rotorB_nxt8(rotorB_mode[8]),
    .rotorB_nxt9(rotorB_mode[9]),
    .rotorB_nxt10(rotorB_mode[10]),
    .rotorB_nxt11(rotorB_mode[11]),
    .rotorB_nxt12(rotorB_mode[12]),
    .rotorB_nxt13(rotorB_mode[13]),
    .rotorB_nxt14(rotorB_mode[14]),
    .rotorB_nxt15(rotorB_mode[15]),
    .rotorB_nxt16(rotorB_mode[16]),
    .rotorB_nxt17(rotorB_mode[17]),
    .rotorB_nxt18(rotorB_mode[18]),
    .rotorB_nxt19(rotorB_mode[19]),
    .rotorB_nxt20(rotorB_mode[20]),
    .rotorB_nxt21(rotorB_mode[21]),
    .rotorB_nxt22(rotorB_mode[22]),
    .rotorB_nxt23(rotorB_mode[23]),
    .rotorB_nxt24(rotorB_mode[24]),
    .rotorB_nxt25(rotorB_mode[25]),
    .rotorB_nxt26(rotorB_mode[26]),
    .rotorB_nxt27(rotorB_mode[27]),
    .rotorB_nxt28(rotorB_mode[28]),
    .rotorB_nxt29(rotorB_mode[29]),
    .rotorB_nxt30(rotorB_mode[30]),
    .rotorB_nxt31(rotorB_mode[31]),
    .rotorB_nxt32(rotorB_mode[32]),
    .rotorB_nxt33(rotorB_mode[33]),
    .rotorB_nxt34(rotorB_mode[34]),
    .rotorB_nxt35(rotorB_mode[35]),
    .rotorB_nxt36(rotorB_mode[36]),
    .rotorB_nxt37(rotorB_mode[37]),
    .rotorB_nxt38(rotorB_mode[38]),
    .rotorB_nxt39(rotorB_mode[39]),
    .rotorB_nxt40(rotorB_mode[40]),
    .rotorB_nxt41(rotorB_mode[41]),
    .rotorB_nxt42(rotorB_mode[42]),
    .rotorB_nxt43(rotorB_mode[43]),
    .rotorB_nxt44(rotorB_mode[44]),
    .rotorB_nxt45(rotorB_mode[45]),
    .rotorB_nxt46(rotorB_mode[46]),
    .rotorB_nxt47(rotorB_mode[47]),
    .rotorB_nxt48(rotorB_mode[48]),
    .rotorB_nxt49(rotorB_mode[49]),
    .rotorB_nxt50(rotorB_mode[50]),
    .rotorB_nxt51(rotorB_mode[51]),
    .rotorB_nxt52(rotorB_mode[52]),
    .rotorB_nxt53(rotorB_mode[53]),
    .rotorB_nxt54(rotorB_mode[54]),
    .rotorB_nxt55(rotorB_mode[55]),
    .rotorB_nxt56(rotorB_mode[56]),
    .rotorB_nxt57(rotorB_mode[57]),
    .rotorB_nxt58(rotorB_mode[58]),
    .rotorB_nxt59(rotorB_mode[59]),
    .rotorB_nxt60(rotorB_mode[60]),
    .rotorB_nxt61(rotorB_mode[61]),
    .rotorB_nxt62(rotorB_mode[62]),
    .rotorB_nxt63(rotorB_mode[63]),
	.rotorB0(rotorB[0]),
    .rotorB1(rotorB[1]),
    .rotorB2(rotorB[2]),
    .rotorB3(rotorB[3]),
    .rotorB4(rotorB[4]),
    .rotorB5(rotorB[5]),
    .rotorB6(rotorB[6]),
    .rotorB7(rotorB[7]),
    .rotorB8(rotorB[8]),
    .rotorB9(rotorB[9]),
    .rotorB10(rotorB[10]),
    .rotorB11(rotorB[11]),
    .rotorB12(rotorB[12]),
    .rotorB13(rotorB[13]),
    .rotorB14(rotorB[14]),
    .rotorB15(rotorB[15]),
    .rotorB16(rotorB[16]),
    .rotorB17(rotorB[17]),
    .rotorB18(rotorB[18]),
    .rotorB19(rotorB[19]),
    .rotorB20(rotorB[20]),
    .rotorB21(rotorB[21]),
    .rotorB22(rotorB[22]),
    .rotorB23(rotorB[23]),
    .rotorB24(rotorB[24]),
    .rotorB25(rotorB[25]),
    .rotorB26(rotorB[26]),
    .rotorB27(rotorB[27]),
    .rotorB28(rotorB[28]),
    .rotorB29(rotorB[29]),
    .rotorB30(rotorB[30]),
    .rotorB31(rotorB[31]),
    .rotorB32(rotorB[32]),
    .rotorB33(rotorB[33]),
    .rotorB34(rotorB[34]),
    .rotorB35(rotorB[35]),
    .rotorB36(rotorB[36]),
    .rotorB37(rotorB[37]),
    .rotorB38(rotorB[38]),
    .rotorB39(rotorB[39]),
    .rotorB40(rotorB[40]),
    .rotorB41(rotorB[41]),
    .rotorB42(rotorB[42]),
    .rotorB43(rotorB[43]),
    .rotorB44(rotorB[44]),
    .rotorB45(rotorB[45]),
    .rotorB46(rotorB[46]),
    .rotorB47(rotorB[47]),
    .rotorB48(rotorB[48]),
    .rotorB49(rotorB[49]),
    .rotorB50(rotorB[50]),
    .rotorB51(rotorB[51]),
    .rotorB52(rotorB[52]),
    .rotorB53(rotorB[53]),
    .rotorB54(rotorB[54]),
    .rotorB55(rotorB[55]),
    .rotorB56(rotorB[56]),
    .rotorB57(rotorB[57]),
    .rotorB58(rotorB[58]),
    .rotorB59(rotorB[59]),
    .rotorB60(rotorB[60]),
    .rotorB61(rotorB[61]),
    .rotorB62(rotorB[62]),
    .rotorB63(rotorB[63])
);

plugboard p(
	.clk(clk),
	.table_idx_buf(table_idx_buf),
	.load_buf(load_buf),
	.code_in_buf(code_in_buf),
	.plugboard0(plugboard[0]),
    .plugboard1(plugboard[1]),
    .plugboard2(plugboard[2]),
    .plugboard3(plugboard[3]),
    .plugboard4(plugboard[4]),
    .plugboard5(plugboard[5]),
    .plugboard6(plugboard[6]),
    .plugboard7(plugboard[7]),
    .plugboard8(plugboard[8]),
    .plugboard9(plugboard[9]),
    .plugboard10(plugboard[10]),
    .plugboard11(plugboard[11]),
    .plugboard12(plugboard[12]),
    .plugboard13(plugboard[13]),
    .plugboard14(plugboard[14]),
    .plugboard15(plugboard[15]),
    .plugboard16(plugboard[16]),
    .plugboard17(plugboard[17]),
    .plugboard18(plugboard[18]),
    .plugboard19(plugboard[19]),
    .plugboard20(plugboard[20]),
    .plugboard21(plugboard[21]),
    .plugboard22(plugboard[22]),
    .plugboard23(plugboard[23]),
    .plugboard24(plugboard[24]),
    .plugboard25(plugboard[25]),
    .plugboard26(plugboard[26]),
    .plugboard27(plugboard[27]),
    .plugboard28(plugboard[28]),
    .plugboard29(plugboard[29]),
    .plugboard30(plugboard[30]),
    .plugboard31(plugboard[31])
);

shift s(
    .clk(clk),
    .crypt_mode_buf(crypt_mode_buf),
    .encrypt_buf(encrypt_buf),
    .encrypt_pipe(encrypt_pipe),
    .rotorA_forward(rotorA_forward[5:4]),
    .rotorB_backward_pipe(rotorB_backward_pipe[5:4]),
    .shift_backward(shift_backward),
    .shift_accu(shift_accu),
    .shift_accu_pipe(shift_accu_pipe)
);

rotorA_forward forward_a(
	.encrypt_pipe(encrypt_pipe), 
	.crypt_mode_buf(crypt_mode_buf), 
	.code_in_1(code_in_1), 
	.code_in_2(code_in_2),
	.code_in_3(code_in_3),
	.out(rotorA_forward)
);

rotorB_forward forward_b(
	.rotorA_forward(rotorA_forward),
	.rotorB0(rotorB[0]),
    .rotorB1(rotorB[1]),
    .rotorB2(rotorB[2]),
    .rotorB3(rotorB[3]),
    .rotorB4(rotorB[4]),
    .rotorB5(rotorB[5]),
    .rotorB6(rotorB[6]),
    .rotorB7(rotorB[7]),
    .rotorB8(rotorB[8]),
    .rotorB9(rotorB[9]),
    .rotorB10(rotorB[10]),
    .rotorB11(rotorB[11]),
    .rotorB12(rotorB[12]),
    .rotorB13(rotorB[13]),
    .rotorB14(rotorB[14]),
    .rotorB15(rotorB[15]),
    .rotorB16(rotorB[16]),
    .rotorB17(rotorB[17]),
    .rotorB18(rotorB[18]),
    .rotorB19(rotorB[19]),
    .rotorB20(rotorB[20]),
    .rotorB21(rotorB[21]),
    .rotorB22(rotorB[22]),
    .rotorB23(rotorB[23]),
    .rotorB24(rotorB[24]),
    .rotorB25(rotorB[25]),
    .rotorB26(rotorB[26]),
    .rotorB27(rotorB[27]),
    .rotorB28(rotorB[28]),
    .rotorB29(rotorB[29]),
    .rotorB30(rotorB[30]),
    .rotorB31(rotorB[31]),
    .rotorB32(rotorB[32]),
    .rotorB33(rotorB[33]),
    .rotorB34(rotorB[34]),
    .rotorB35(rotorB[35]),
    .rotorB36(rotorB[36]),
    .rotorB37(rotorB[37]),
    .rotorB38(rotorB[38]),
    .rotorB39(rotorB[39]),
    .rotorB40(rotorB[40]),
    .rotorB41(rotorB[41]),
    .rotorB42(rotorB[42]),
    .rotorB43(rotorB[43]),
    .rotorB44(rotorB[44]),
    .rotorB45(rotorB[45]),
    .rotorB46(rotorB[46]),
    .rotorB47(rotorB[47]),
    .rotorB48(rotorB[48]),
    .rotorB49(rotorB[49]),
    .rotorB50(rotorB[50]),
    .rotorB51(rotorB[51]),
    .rotorB52(rotorB[52]),
    .rotorB53(rotorB[53]),
    .rotorB54(rotorB[54]),
    .rotorB55(rotorB[55]),
    .rotorB56(rotorB[56]),
    .rotorB57(rotorB[57]),
    .rotorB58(rotorB[58]),
    .rotorB59(rotorB[59]),
    .rotorB60(rotorB[60]),
    .rotorB61(rotorB[61]),
    .rotorB62(rotorB[62]),
    .rotorB63(rotorB[63]),
	.out(rotorB_forward)
);

plugboard_forward pf(
	.rotorB_forward(rotorB_forward),
	.plugboard0(plugboard[0]),
    .plugboard1(plugboard[1]),
    .plugboard2(plugboard[2]),
    .plugboard3(plugboard[3]),
    .plugboard4(plugboard[4]),
    .plugboard5(plugboard[5]),
    .plugboard6(plugboard[6]),
    .plugboard7(plugboard[7]),
    .plugboard8(plugboard[8]),
    .plugboard9(plugboard[9]),
    .plugboard10(plugboard[10]),
    .plugboard11(plugboard[11]),
    .plugboard12(plugboard[12]),
    .plugboard13(plugboard[13]),
    .plugboard14(plugboard[14]),
    .plugboard15(plugboard[15]),
    .plugboard16(plugboard[16]),
    .plugboard17(plugboard[17]),
    .plugboard18(plugboard[18]),
    .plugboard19(plugboard[19]),
    .plugboard20(plugboard[20]),
    .plugboard21(plugboard[21]),
    .plugboard22(plugboard[22]),
    .plugboard23(plugboard[23]),
    .plugboard24(plugboard[24]),
    .plugboard25(plugboard[25]),
    .plugboard26(plugboard[26]),
    .plugboard27(plugboard[27]),
    .plugboard28(plugboard[28]),
    .plugboard29(plugboard[29]),
    .plugboard30(plugboard[30]),
    .plugboard31(plugboard[31]),
	.out(plugboard_forward)
);

plugboard_backward pb(
	.plugboard_forward(plugboard_forward),
	.plugboard0(plugboard[0]),
    .plugboard1(plugboard[1]),
    .plugboard2(plugboard[2]),
    .plugboard3(plugboard[3]),
    .plugboard4(plugboard[4]),
    .plugboard5(plugboard[5]),
    .plugboard6(plugboard[6]),
    .plugboard7(plugboard[7]),
    .plugboard8(plugboard[8]),
    .plugboard9(plugboard[9]),
    .plugboard10(plugboard[10]),
    .plugboard11(plugboard[11]),
    .plugboard12(plugboard[12]),
    .plugboard13(plugboard[13]),
    .plugboard14(plugboard[14]),
    .plugboard15(plugboard[15]),
    .plugboard16(plugboard[16]),
    .plugboard17(plugboard[17]),
    .plugboard18(plugboard[18]),
    .plugboard19(plugboard[19]),
    .plugboard20(plugboard[20]),
    .plugboard21(plugboard[21]),
    .plugboard22(plugboard[22]),
    .plugboard23(plugboard[23]),
    .plugboard24(plugboard[24]),
    .plugboard25(plugboard[25]),
    .plugboard26(plugboard[26]),
    .plugboard27(plugboard[27]),
    .plugboard28(plugboard[28]),
    .plugboard29(plugboard[29]),
    .plugboard30(plugboard[30]),
    .plugboard31(plugboard[31]),
	.out(plugboard_backward)
);

rotorB_backward backward_b(
	.rotorB0(rotorB[0]),
    .rotorB1(rotorB[1]),
    .rotorB2(rotorB[2]),
    .rotorB3(rotorB[3]),
    .rotorB4(rotorB[4]),
    .rotorB5(rotorB[5]),
    .rotorB6(rotorB[6]),
    .rotorB7(rotorB[7]),
    .rotorB8(rotorB[8]),
    .rotorB9(rotorB[9]),
    .rotorB10(rotorB[10]),
    .rotorB11(rotorB[11]),
    .rotorB12(rotorB[12]),
    .rotorB13(rotorB[13]),
    .rotorB14(rotorB[14]),
    .rotorB15(rotorB[15]),
    .rotorB16(rotorB[16]),
    .rotorB17(rotorB[17]),
    .rotorB18(rotorB[18]),
    .rotorB19(rotorB[19]),
    .rotorB20(rotorB[20]),
    .rotorB21(rotorB[21]),
    .rotorB22(rotorB[22]),
    .rotorB23(rotorB[23]),
    .rotorB24(rotorB[24]),
    .rotorB25(rotorB[25]),
    .rotorB26(rotorB[26]),
    .rotorB27(rotorB[27]),
    .rotorB28(rotorB[28]),
    .rotorB29(rotorB[29]),
    .rotorB30(rotorB[30]),
    .rotorB31(rotorB[31]),
    .rotorB32(rotorB[32]),
    .rotorB33(rotorB[33]),
    .rotorB34(rotorB[34]),
    .rotorB35(rotorB[35]),
    .rotorB36(rotorB[36]),
    .rotorB37(rotorB[37]),
    .rotorB38(rotorB[38]),
    .rotorB39(rotorB[39]),
    .rotorB40(rotorB[40]),
    .rotorB41(rotorB[41]),
    .rotorB42(rotorB[42]),
    .rotorB43(rotorB[43]),
    .rotorB44(rotorB[44]),
    .rotorB45(rotorB[45]),
    .rotorB46(rotorB[46]),
    .rotorB47(rotorB[47]),
    .rotorB48(rotorB[48]),
    .rotorB49(rotorB[49]),
    .rotorB50(rotorB[50]),
    .rotorB51(rotorB[51]),
    .rotorB52(rotorB[52]),
    .rotorB53(rotorB[53]),
    .rotorB54(rotorB[54]),
    .rotorB55(rotorB[55]),
    .rotorB56(rotorB[56]),
    .rotorB57(rotorB[57]),
    .rotorB58(rotorB[58]),
    .rotorB59(rotorB[59]),
    .rotorB60(rotorB[60]),
    .rotorB61(rotorB[61]),
    .rotorB62(rotorB[62]),
    .rotorB63(rotorB[63]),
	.plugboard_backward(plugboard_backward),
	.out(rotorB_backward)
);

rotorA_backward backward_a(
	.crypt_mode_buf(crypt_mode_buf),
	.rotorA0(rotorA[0]),
    .rotorA1(rotorA[1]),
    .rotorA2(rotorA[2]),
    .rotorA3(rotorA[3]),
    .rotorA4(rotorA[4]),
    .rotorA5(rotorA[5]),
    .rotorA6(rotorA[6]),
    .rotorA7(rotorA[7]),
    .rotorA8(rotorA[8]),
    .rotorA9(rotorA[9]),
    .rotorA10(rotorA[10]),
    .rotorA11(rotorA[11]),
    .rotorA12(rotorA[12]),
    .rotorA13(rotorA[13]),
    .rotorA14(rotorA[14]),
    .rotorA15(rotorA[15]),
    .rotorA16(rotorA[16]),
    .rotorA17(rotorA[17]),
    .rotorA18(rotorA[18]),
    .rotorA19(rotorA[19]),
    .rotorA20(rotorA[20]),
    .rotorA21(rotorA[21]),
    .rotorA22(rotorA[22]),
    .rotorA23(rotorA[23]),
    .rotorA24(rotorA[24]),
    .rotorA25(rotorA[25]),
    .rotorA26(rotorA[26]),
    .rotorA27(rotorA[27]),
    .rotorA28(rotorA[28]),
    .rotorA29(rotorA[29]),
    .rotorA30(rotorA[30]),
    .rotorA31(rotorA[31]),
    .rotorA32(rotorA[32]),
    .rotorA33(rotorA[33]),
    .rotorA34(rotorA[34]),
    .rotorA35(rotorA[35]),
    .rotorA36(rotorA[36]),
    .rotorA37(rotorA[37]),
    .rotorA38(rotorA[38]),
    .rotorA39(rotorA[39]),
    .rotorA40(rotorA[40]),
    .rotorA41(rotorA[41]),
    .rotorA42(rotorA[42]),
    .rotorA43(rotorA[43]),
    .rotorA44(rotorA[44]),
    .rotorA45(rotorA[45]),
    .rotorA46(rotorA[46]),
    .rotorA47(rotorA[47]),
    .rotorA48(rotorA[48]),
    .rotorA49(rotorA[49]),
    .rotorA50(rotorA[50]),
    .rotorA51(rotorA[51]),
    .rotorA52(rotorA[52]),
    .rotorA53(rotorA[53]),
    .rotorA54(rotorA[54]),
    .rotorA55(rotorA[55]),
    .rotorA56(rotorA[56]),
    .rotorA57(rotorA[57]),
    .rotorA58(rotorA[58]),
    .rotorA59(rotorA[59]),
    .rotorA60(rotorA[60]),
    .rotorA61(rotorA[61]),
    .rotorA62(rotorA[62]),
    .rotorA63(rotorA[63]),
	.rotorB_backward_pipe(rotorB_backward_pipe),
	.shift_accu(shift_accu),
	.shift_accu_pipe(shift_accu_pipe),
	.out(code_out_nxt)
);

mode m(
	.encrypt_buf(encrypt_buf),
	.crypt_mode_buf(crypt_mode_buf),
	.plugboard_backward(plugboard_backward[1:0]),
	.rotorB_forward(rotorB_forward[1:0]),
	.rotorB0(rotorB[0]),
    .rotorB1(rotorB[1]),
    .rotorB2(rotorB[2]),
    .rotorB3(rotorB[3]),
    .rotorB4(rotorB[4]),
    .rotorB5(rotorB[5]),
    .rotorB6(rotorB[6]),
    .rotorB7(rotorB[7]),
    .rotorB8(rotorB[8]),
    .rotorB9(rotorB[9]),
    .rotorB10(rotorB[10]),
    .rotorB11(rotorB[11]),
    .rotorB12(rotorB[12]),
    .rotorB13(rotorB[13]),
    .rotorB14(rotorB[14]),
    .rotorB15(rotorB[15]),
    .rotorB16(rotorB[16]),
    .rotorB17(rotorB[17]),
    .rotorB18(rotorB[18]),
    .rotorB19(rotorB[19]),
    .rotorB20(rotorB[20]),
    .rotorB21(rotorB[21]),
    .rotorB22(rotorB[22]),
    .rotorB23(rotorB[23]),
    .rotorB24(rotorB[24]),
    .rotorB25(rotorB[25]),
    .rotorB26(rotorB[26]),
    .rotorB27(rotorB[27]),
    .rotorB28(rotorB[28]),
    .rotorB29(rotorB[29]),
    .rotorB30(rotorB[30]),
    .rotorB31(rotorB[31]),
    .rotorB32(rotorB[32]),
    .rotorB33(rotorB[33]),
    .rotorB34(rotorB[34]),
    .rotorB35(rotorB[35]),
    .rotorB36(rotorB[36]),
    .rotorB37(rotorB[37]),
    .rotorB38(rotorB[38]),
    .rotorB39(rotorB[39]),
    .rotorB40(rotorB[40]),
    .rotorB41(rotorB[41]),
    .rotorB42(rotorB[42]),
    .rotorB43(rotorB[43]),
    .rotorB44(rotorB[44]),
    .rotorB45(rotorB[45]),
    .rotorB46(rotorB[46]),
    .rotorB47(rotorB[47]),
    .rotorB48(rotorB[48]),
    .rotorB49(rotorB[49]),
    .rotorB50(rotorB[50]),
    .rotorB51(rotorB[51]),
    .rotorB52(rotorB[52]),
    .rotorB53(rotorB[53]),
    .rotorB54(rotorB[54]),
    .rotorB55(rotorB[55]),
    .rotorB56(rotorB[56]),
    .rotorB57(rotorB[57]),
    .rotorB58(rotorB[58]),
    .rotorB59(rotorB[59]),
    .rotorB60(rotorB[60]),
    .rotorB61(rotorB[61]),
    .rotorB62(rotorB[62]),
    .rotorB63(rotorB[63]),
	.rotorB_nxt0(rotorB_mode[0]),
    .rotorB_nxt1(rotorB_mode[1]),
    .rotorB_nxt2(rotorB_mode[2]),
    .rotorB_nxt3(rotorB_mode[3]),
    .rotorB_nxt4(rotorB_mode[4]),
    .rotorB_nxt5(rotorB_mode[5]),
    .rotorB_nxt6(rotorB_mode[6]),
    .rotorB_nxt7(rotorB_mode[7]),
    .rotorB_nxt8(rotorB_mode[8]),
    .rotorB_nxt9(rotorB_mode[9]),
    .rotorB_nxt10(rotorB_mode[10]),
    .rotorB_nxt11(rotorB_mode[11]),
    .rotorB_nxt12(rotorB_mode[12]),
    .rotorB_nxt13(rotorB_mode[13]),
    .rotorB_nxt14(rotorB_mode[14]),
    .rotorB_nxt15(rotorB_mode[15]),
    .rotorB_nxt16(rotorB_mode[16]),
    .rotorB_nxt17(rotorB_mode[17]),
    .rotorB_nxt18(rotorB_mode[18]),
    .rotorB_nxt19(rotorB_mode[19]),
    .rotorB_nxt20(rotorB_mode[20]),
    .rotorB_nxt21(rotorB_mode[21]),
    .rotorB_nxt22(rotorB_mode[22]),
    .rotorB_nxt23(rotorB_mode[23]),
    .rotorB_nxt24(rotorB_mode[24]),
    .rotorB_nxt25(rotorB_mode[25]),
    .rotorB_nxt26(rotorB_mode[26]),
    .rotorB_nxt27(rotorB_mode[27]),
    .rotorB_nxt28(rotorB_mode[28]),
    .rotorB_nxt29(rotorB_mode[29]),
    .rotorB_nxt30(rotorB_mode[30]),
    .rotorB_nxt31(rotorB_mode[31]),
    .rotorB_nxt32(rotorB_mode[32]),
    .rotorB_nxt33(rotorB_mode[33]),
    .rotorB_nxt34(rotorB_mode[34]),
    .rotorB_nxt35(rotorB_mode[35]),
    .rotorB_nxt36(rotorB_mode[36]),
    .rotorB_nxt37(rotorB_mode[37]),
    .rotorB_nxt38(rotorB_mode[38]),
    .rotorB_nxt39(rotorB_mode[39]),
    .rotorB_nxt40(rotorB_mode[40]),
    .rotorB_nxt41(rotorB_mode[41]),
    .rotorB_nxt42(rotorB_mode[42]),
    .rotorB_nxt43(rotorB_mode[43]),
    .rotorB_nxt44(rotorB_mode[44]),
    .rotorB_nxt45(rotorB_mode[45]),
    .rotorB_nxt46(rotorB_mode[46]),
    .rotorB_nxt47(rotorB_mode[47]),
    .rotorB_nxt48(rotorB_mode[48]),
    .rotorB_nxt49(rotorB_mode[49]),
    .rotorB_nxt50(rotorB_mode[50]),
    .rotorB_nxt51(rotorB_mode[51]),
    .rotorB_nxt52(rotorB_mode[52]),
    .rotorB_nxt53(rotorB_mode[53]),
    .rotorB_nxt54(rotorB_mode[54]),
    .rotorB_nxt55(rotorB_mode[55]),
    .rotorB_nxt56(rotorB_mode[56]),
    .rotorB_nxt57(rotorB_mode[57]),
    .rotorB_nxt58(rotorB_mode[58]),
    .rotorB_nxt59(rotorB_mode[59]),
    .rotorB_nxt60(rotorB_mode[60]),
    .rotorB_nxt61(rotorB_mode[61]),
    .rotorB_nxt62(rotorB_mode[62]),
    .rotorB_nxt63(rotorB_mode[63])
);

endmodule